module cla_4(
  input 
);
    
endmodule //cla_4
